//--------------------------------------------------------------
//  dispatcher.v
//  -----------------------------------------------------------
//  1. 功能 : 從佇列 FIFO 取出一筆資料，依序派發給
//            第一個「空閒」的櫃檯 (counter)。
//  2. 規則 : 固定優先權  櫃檯1 → 櫃檯2 → 櫃檯3
//            只要成功派發，就對 FIFO 送出 re=1 讀脈衝。
//  3. 時序 : 以 clk 正緣為基準，所有旗標皆同步重設。
//--------------------------------------------------------------
module dispatcher(clk, rst_n, empty, busy, qn, qt, re, ld, dn, dt);
    parameter DT_SZ = 4;        // 資料大小，預設 4 bits
    parameter CNTER = 3;        // 櫃台數量
	//==================== 時脈 / 重設 =========================
    input  clk;
    input  rst_n;               // 同步低有效

    //==================== 來自 FIFO 的訊號 ====================
    input        empty;         // =1 代表 FIFO 為空
    input  [DT_SZ-1:0] qn;      // 佇列首端客人編號
    input  [DT_SZ-1:0] qt;      // 佇列首端服務時間

    //==================== 各櫃檯忙碌狀態 ======================
    // busy[i] = 1  該櫃檯正在服務，不可派發
    input  [CNTER-1:0] busy;

    //==================== 給 FIFO 的控制 ======================
    output reg   re;            // 讀出脈衝 (HIGH 1 個 clk)

    //==================== 給三個 counter 的載入控制 ===========
    // ld?  : 載入脈衝 (HIGH 1 個 clk)
    // dn?/dt? : 欲載入之 {編號, 時間}
    output reg [CNTER-1:0] ld;
	output reg [DT_SZ-1:0] dn;
	output reg [DT_SZ-1:0] dt;

	// for 迴圈用
	integer i;

	//--------------------------------------------------------------
	//  派發邏輯
	//--------------------------------------------------------------
	always @(posedge clk or negedge rst_n) begin
		if (!rst_n) begin
			// --------- 非同步重設 ---------------------------------
			re  <= 1'b0;
			ld <= {CNTER{1'b0}}; // 脈衝清 0
			dn <= {DT_SZ{1'b0}}; // 暫存清 0
			dt <= {DT_SZ{1'b0}}; // 暫存清 0
		end
		else begin
			#2
			// --------- 預設值：每拍先清脈衝 ----------------------------
			re  <= 1'b0;
			ld <= {CNTER{1'b0}};      // 脈衝清 0
			// --------- 當 FIFO 非空，嘗試派發 ----------------------
			if (!empty) begin:block
				for (i = 0; i < CNTER; i = i + 1) begin
					if (!busy[i]) begin
						re <= 1'b1; 
						ld[i] <= 1'b1;
						dn <= qn;
						dt <= qt;
						disable block; // 找到空位就退出 for 迴圈
					end
				end
				// 若全忙碌：不派發，re=0，資料留在 FIFO
			end
		end
	end
endmodule